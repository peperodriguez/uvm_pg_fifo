module top;
  
  tb t();

endmodule